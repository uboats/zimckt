VDD 103 0 DC 3
Vword 110 0 DC 3
Vbit 120 0 DC 3
Vbitb 130 0 DC 3

vin 102 0 DC 0

*    d     g     s
M1 104 102 103 p 30e-6 0.35e-6 1
M2 104 102 0 n 10e-6 0.35e-6 2

M3 102 104 103 p 30e-6 0.35e-6 1
M4 102 104 0 n 10e-6 0.35e-6 2

Ma 105 110 102 n 10e-6 0.35e-6 2
R1 120 105 10

Mb 108 110 104 n 10e-6 0.35e-6 2
R2 130 108 1000

.MODEL 1 VT -0.75 MU 5e-2 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14
.MODEL 2 VT 0.83 MU 1.5e-1 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14

.DC SWEEP vin 0 3 0.02
*.DC
.PLOTNV 104
.PLOTNV 102
