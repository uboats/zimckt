* ckt file for parser

* interpret this as a voltage step

Vdriver1 256 0 1


* port 256 - load 2.000000e+00

r1	256	261	9.999000e+00
c2	261	0	9.999e-14
r3	261	262	9.999000e+00
c4	262	0	9.999e-14
r5	262	129	9.999000e+00

r6	129	263	2.381700e+01
c7	263	0	2.3817e-13
r8	263	264	2.381700e+01
c9	264	0	2.3817e-13
r10	264	130	2.381700e+01

r11	129	265	2.381800e+01
c12	265	0	2.3818e-13
r13	265	266	2.381800e+01
c14	266	0	2.3818e-13
r15	266	131	2.381800e+01

r16	130	267	1.622400e+01
c17	267	0	1.6224e-13
r18	267	268	1.622400e+01
c19	268	0	1.6224e-13
r20	268	132	1.622400e+01

r21	130	269	1.622300e+01
c22	269	0	1.6223e-13
r23	269	270	1.622300e+01
c24	270	0	1.6223e-13
r25	270	133	1.622300e+01

r26	131	271	1.147100e+01
c27	271	0	1.1471e-13
r28	271	272	1.147100e+01
c29	272	0	1.1471e-13
r30	272	134	1.147100e+01

r31	131	273	1.147200e+01
c32	273	0	1.1472e-13
r33	273	274	1.147200e+01
c34	274	0	1.1472e-13
r35	274	135	1.147200e+01

r36	132	275	1.173700e+01
c37	275	0	1.1737e-13
r38	275	276	1.173700e+01
c39	276	0	1.1737e-13
r40	276	136	1.173700e+01

r41	132	277	1.173700e+01
c42	277	0	1.1737e-13
r43	277	278	1.173700e+01
c44	278	0	1.1737e-13
r45	278	137	1.173700e+01

r46	136	279	1.050100e+01
c47	279	0	1.0501e-13
r48	279	280	1.050100e+01
c49	280	0	1.0501e-13
r50	280	138	1.050100e+01

r51	136	281	1.050000e+01
c52	281	0	1.05e-13
r53	281	282	1.050000e+01
c54	282	0	1.05e-13
r55	282	139	1.050000e+01

r56	137	283	7.556000e+00
c57	283	0	7.556e-14
r58	283	284	7.556000e+00
c59	284	0	7.556e-14
r60	284	140	7.556000e+00

r61	137	285	7.555000e+00
c62	285	0	7.555e-14
r63	285	286	7.555000e+00
c64	286	0	7.555e-14
r65	286	141	7.555000e+00

r66	138	287	7.719000e+00
c67	287	0	7.719e-14
r68	287	288	7.719000e+00
c69	288	0	7.719e-14
r70	288	142	7.719000e+00

r71	138	289	7.720000e+00
c72	289	0	7.72e-14
r73	289	290	7.720000e+00
c74	290	0	7.72e-14
r75	290	143	7.720000e+00

r76	142	291	7.666000e+00
c77	291	0	7.666e-14
r78	291	292	7.666000e+00
c79	292	0	7.666e-14
r80	292	144	7.666000e+00

r81	142	293	7.666000e+00
c82	293	0	7.666e-14
r83	293	294	7.666000e+00
c84	294	0	7.666e-14
r85	294	145	7.666000e+00

r86	143	295	1.161500e+01
c87	295	0	1.1615e-13
r88	295	296	1.161500e+01
c89	296	0	1.1615e-13
r90	296	146	1.161500e+01

r91	143	297	1.161500e+01
c92	297	0	1.1615e-13
r93	297	298	1.161500e+01
c94	298	0	1.1615e-13
r95	298	147	1.161500e+01

r96	144	299	6.494000e+00
c97	299	0	6.494e-14
r98	299	300	6.494000e+00
c99	300	0	6.494e-14
r100	300	41	6.494000e+00

* port 41 - load 3.100000e-02

r101	144	301	6.494000e+00
c102	301	0	6.494e-14
r103	301	302	6.494000e+00
c104	302	0	6.494e-14
r105	302	42	6.494000e+00

* port 42 - load 7.500000e-02

r106	145	303	8.438000e+00
c107	303	0	8.438e-14
r108	303	304	8.438000e+00
c109	304	0	8.438e-14
r110	304	82	8.438000e+00

* port 82 - load 4.900000e-02

r111	145	305	8.438000e+00
c112	305	0	8.438e-14
r113	305	306	8.438000e+00
c114	306	0	8.438e-14
r115	306	40	8.438000e+00

* port 40 - load 5.300000e-02

r116	146	307	8.330000e+00
c117	307	0	8.33e-14
r118	307	308	8.330000e+00
c119	308	0	8.33e-14
r120	308	43	8.330000e+00

* port 43 - load 3.400000e-02

r121	146	309	8.330000e+00
c122	309	0	8.33e-14
r123	309	310	8.330000e+00
c124	310	0	8.33e-14
r125	310	48	8.330000e+00

* port 48 - load 7.800000e-02

r126	147	311	5.940000e-01
c127	311	0	5.94e-15
r128	311	312	5.940000e-01
c129	312	0	5.94e-15
r130	312	85	5.940000e-01

* port 85 - load 7.800000e-02

r131	147	313	5.930000e-01
c132	313	0	5.93e-15
r133	313	314	5.930000e-01
c134	314	0	5.93e-15
r135	314	50	5.930000e-01

* port 50 - load 4.200000e-02

r136	139	315	5.136000e+00
c137	315	0	5.136e-14
r138	315	316	5.136000e+00
c139	316	0	5.136e-14
r140	316	148	5.136000e+00

r141	139	317	5.137000e+00
c142	317	0	5.137e-14
r143	317	318	5.137000e+00
c144	318	0	5.137e-14
r145	318	149	5.137000e+00

r146	148	319	5.351000e+00
c147	319	0	5.351e-14
r148	319	320	5.351000e+00
c149	320	0	5.351e-14
r150	320	150	5.351000e+00

r151	148	321	5.351000e+00
c152	321	0	5.351e-14
r153	321	322	5.351000e+00
c154	322	0	5.351e-14
r155	322	151	5.351000e+00

r156	149	323	2.714000e+00
c157	323	0	2.714e-14
r158	323	324	2.714000e+00
c159	324	0	2.714e-14
r160	324	152	2.714000e+00

r161	149	325	2.714000e+00
c162	325	0	2.714e-14
r163	325	326	2.714000e+00
c164	326	0	2.714e-14
r165	326	153	2.714000e+00

r166	150	327	3.408000e+00
c167	327	0	3.408e-14
r168	327	328	3.408000e+00
c169	328	0	3.408e-14
r170	328	83	3.408000e+00

* port 83 - load 3.100000e-02

r171	150	329	3.409000e+00
c172	329	0	3.409e-14
r173	329	330	3.409000e+00
c174	330	0	3.409e-14
r175	330	81	3.409000e+00

* port 81 - load 6.600000e-02

r176	151	331	1.613000e+00
c177	331	0	1.613e-14
r178	331	332	1.613000e+00
c179	332	0	1.613e-14
r180	332	77	1.613000e+00

* port 77 - load 7.900000e-02

r181	151	333	1.613000e+00
c182	333	0	1.613e-14
r183	333	334	1.613000e+00
c184	334	0	1.613e-14
r185	334	84	1.613000e+00

* port 84 - load 6.400000e-02

r186	152	335	4.870000e-01
c187	335	0	4.87e-15
r188	335	336	4.870000e-01
c189	336	0	4.87e-15
r190	336	80	4.870000e-01

* port 80 - load 3.500000e-02

r191	152	337	4.880000e-01
c192	337	0	4.88e-15
r193	337	338	4.880000e-01
c194	338	0	4.88e-15
r195	338	54	4.880000e-01

* port 54 - load 6.000000e-02

r196	153	339	9.350000e-01
c197	339	0	9.35e-15
r198	339	340	9.350000e-01
c199	340	0	9.35e-15
r200	340	53	9.350000e-01

* port 53 - load 3.300000e-02

r201	153	341	9.350000e-01
c202	341	0	9.35e-15
r203	341	342	9.350000e-01
c204	342	0	9.35e-15
r205	342	51	9.350000e-01

* port 51 - load 4.700000e-02

r206	140	343	5.183000e+00
c207	343	0	5.183e-14
r208	343	344	5.183000e+00
c209	344	0	5.183e-14
r210	344	154	5.183000e+00

r211	140	345	5.183000e+00
c212	345	0	5.183e-14
r213	345	346	5.183000e+00
c214	346	0	5.183e-14
r215	346	155	5.183000e+00

r216	154	347	6.147000e+00
c217	347	0	6.147e-14
r218	347	348	6.147000e+00
c219	348	0	6.147e-14
r220	348	156	6.147000e+00

r221	154	349	6.145000e+00
c222	349	0	6.145e-14
r223	349	350	6.145000e+00
c224	350	0	6.145e-14
r225	350	157	6.145000e+00

r226	155	351	2.516000e+00
c227	351	0	2.516e-14
r228	351	352	2.516000e+00
c229	352	0	2.516e-14
r230	352	158	2.516000e+00

r231	155	353	2.516000e+00
c232	353	0	2.516e-14
r233	353	354	2.516000e+00
c234	354	0	2.516e-14
r235	354	159	2.516000e+00

r236	156	355	2.475000e+00
c237	355	0	2.475e-14
r238	355	356	2.475000e+00
c239	356	0	2.475e-14
r240	356	38	2.475000e+00

* port 38 - load 6.700000e-02

r241	156	357	2.474000e+00
c242	357	0	2.474e-14
r243	357	358	2.474000e+00
c244	358	0	2.474e-14
r245	358	44	2.474000e+00

* port 44 - load 6.300000e-02

r246	157	359	3.420000e+00
c247	359	0	3.42e-14
r248	359	360	3.420000e+00
c249	360	0	3.42e-14
r250	360	39	3.420000e+00

* port 39 - load 3.500000e-02

r251	157	361	3.419000e+00
c252	361	0	3.419e-14
r253	361	362	3.419000e+00
c254	362	0	3.419e-14
r255	362	47	3.419000e+00

* port 47 - load 7.000000e-02

r256	158	363	3.997000e+00
c257	363	0	3.997e-14
r258	363	364	3.997000e+00
c259	364	0	3.997e-14
r260	364	45	3.997000e+00

* port 45 - load 4.500000e-02

r261	158	365	3.998000e+00
c262	365	0	3.998e-14
r263	365	366	3.998000e+00
c264	366	0	3.998e-14
r265	366	37	3.998000e+00

* port 37 - load 8.000000e-02

r266	159	367	3.160000e-01
c267	367	0	3.16e-15
r268	367	368	3.160000e-01
c269	368	0	3.16e-15
r270	368	36	3.160000e-01

* port 36 - load 6.300000e-02

r271	159	369	3.170000e-01
c272	369	0	3.17e-15
r273	369	370	3.170000e-01
c274	370	0	3.17e-15
r275	370	89	3.170000e-01

* port 89 - load 5.800000e-02

r276	141	371	2.802000e+00
c277	371	0	2.802e-14
r278	371	372	2.802000e+00
c279	372	0	2.802e-14
r280	372	160	2.802000e+00

r281	141	373	2.801000e+00
c282	373	0	2.801e-14
r283	373	374	2.801000e+00
c284	374	0	2.801e-14
r285	374	161	2.801000e+00

r286	160	375	5.530000e+00
c287	375	0	5.53e-14
r288	375	376	5.530000e+00
c289	376	0	5.53e-14
r290	376	162	5.530000e+00

r291	160	377	5.532000e+00
c292	377	0	5.532e-14
r293	377	378	5.532000e+00
c294	378	0	5.532e-14
r295	378	163	5.532000e+00

r296	161	379	3.809000e+00
c297	379	0	3.809e-14
r298	379	380	3.809000e+00
c299	380	0	3.809e-14
r300	380	164	3.809000e+00

r301	161	381	3.807000e+00
c302	381	0	3.807e-14
r303	381	382	3.807000e+00
c304	382	0	3.807e-14
r305	382	165	3.807000e+00

r306	162	383	3.628000e+00
c307	383	0	3.628e-14
r308	383	384	3.628000e+00
c309	384	0	3.628e-14
r310	384	49	3.628000e+00

* port 49 - load 7.700000e-02

r311	162	385	3.628000e+00
c312	385	0	3.628e-14
r313	385	386	3.628000e+00
c314	386	0	3.628e-14
r315	386	46	3.628000e+00

* port 46 - load 4.600000e-02

r316	163	387	6.398000e+00
c317	387	0	6.398e-14
r318	387	388	6.398000e+00
c319	388	0	6.398e-14
r320	388	86	6.398000e+00

* port 86 - load 3.400000e-02

r321	163	389	6.399000e+00
c322	389	0	6.399e-14
r323	389	390	6.399000e+00
c324	390	0	6.399e-14
r325	390	1	6.399000e+00

* port 1 - load 5.900000e-02

r326	164	391	2.034000e+00
c327	391	0	2.034e-14
r328	391	392	2.034000e+00
c329	392	0	2.034e-14
r330	392	27	2.034000e+00

* port 27 - load 5.800000e-02

r331	164	393	2.035000e+00
c332	393	0	2.035e-14
r333	393	394	2.035000e+00
c334	394	0	2.035e-14
r335	394	26	2.035000e+00

* port 26 - load 4.100000e-02

r336	165	395	2.737000e+00
c337	395	0	2.737e-14
r338	395	396	2.737000e+00
c339	396	0	2.737e-14
r340	396	87	2.737000e+00

* port 87 - load 4.200000e-02

r341	165	397	2.736000e+00
c342	397	0	2.736e-14
r343	397	398	2.736000e+00
c344	398	0	2.736e-14
r345	398	88	2.736000e+00

* port 88 - load 3.300000e-02

r346	133	399	7.753000e+00
c347	399	0	7.753e-14
r348	399	400	7.753000e+00
c349	400	0	7.753e-14
r350	400	166	7.753000e+00

r351	133	401	7.752000e+00
c352	401	0	7.752e-14
r353	401	402	7.752000e+00
c354	402	0	7.752e-14
r355	402	167	7.752000e+00

r356	166	403	7.848000e+00
c357	403	0	7.848e-14
r358	403	404	7.848000e+00
c359	404	0	7.848e-14
r360	404	168	7.848000e+00

r361	166	405	7.849000e+00
c362	405	0	7.849e-14
r363	405	406	7.849000e+00
c364	406	0	7.849e-14
r365	406	169	7.849000e+00

r366	167	407	3.966000e+00
c367	407	0	3.966e-14
r368	407	408	3.966000e+00
c369	408	0	3.966e-14
r370	408	170	3.966000e+00

r371	167	409	3.966000e+00
c372	409	0	3.966e-14
r373	409	410	3.966000e+00
c374	410	0	3.966e-14
r375	410	171	3.966000e+00

r376	168	411	4.735000e+00
c377	411	0	4.735e-14
r378	411	412	4.735000e+00
c379	412	0	4.735e-14
r380	412	172	4.735000e+00

r381	168	413	4.736000e+00
c382	413	0	4.736e-14
r383	413	414	4.736000e+00
c384	414	0	4.736e-14
r385	414	173	4.736000e+00

r386	172	415	1.158000e+00
c387	415	0	1.158e-14
r388	415	416	1.158000e+00
c389	416	0	1.158e-14
r390	416	174	1.158000e+00

r391	172	417	1.159000e+00
c392	417	0	1.159e-14
r393	417	418	1.159000e+00
c394	418	0	1.159e-14
r395	418	175	1.159000e+00

r396	173	419	2.340000e+00
c397	419	0	2.34e-14
r398	419	420	2.340000e+00
c399	420	0	2.34e-14
r400	420	176	2.340000e+00

r401	173	421	2.341000e+00
c402	421	0	2.341e-14
r403	421	422	2.341000e+00
c404	422	0	2.341e-14
r405	422	177	2.341000e+00

r406	174	423	4.610000e-01
c407	423	0	4.61e-15
r408	423	424	4.610000e-01
c409	424	0	4.61e-15
r410	424	56	4.610000e-01

* port 56 - load 3.900000e-02

r411	174	425	4.610000e-01
c412	425	0	4.61e-15
r413	425	426	4.610000e-01
c414	426	0	4.61e-15
r415	426	55	4.610000e-01

* port 55 - load 4.200000e-02

r416	175	427	5.304000e+00
c417	427	0	5.304e-14
r418	427	428	5.304000e+00
c419	428	0	5.304e-14
r420	428	76	5.304000e+00

* port 76 - load 6.400000e-02

r421	175	429	5.304000e+00
c422	429	0	5.304e-14
r423	429	430	5.304000e+00
c424	430	0	5.304e-14
r425	430	78	5.304000e+00

* port 78 - load 7.200000e-02

r426	176	431	2.683000e+00
c427	431	0	2.683e-14
r428	431	432	2.683000e+00
c429	432	0	2.683e-14
r430	432	67	2.683000e+00

* port 67 - load 3.500000e-02

r431	176	433	2.684000e+00
c432	433	0	2.684e-14
r433	433	434	2.684000e+00
c434	434	0	2.684e-14
r435	434	79	2.684000e+00

* port 79 - load 4.100000e-02

r436	177	435	1.802000e+00
c437	435	0	1.802e-14
r438	435	436	1.802000e+00
c439	436	0	1.802e-14
r440	436	65	1.802000e+00

* port 65 - load 7.700000e-02

r441	177	437	1.801000e+00
c442	437	0	1.801e-14
r443	437	438	1.801000e+00
c444	438	0	1.801e-14
r445	438	57	1.801000e+00

* port 57 - load 6.000000e-02

r446	169	439	2.591000e+00
c447	439	0	2.591e-14
r448	439	440	2.591000e+00
c449	440	0	2.591e-14
r450	440	178	2.591000e+00

r451	169	441	2.590000e+00
c452	441	0	2.59e-14
r453	441	442	2.590000e+00
c454	442	0	2.59e-14
r455	442	179	2.590000e+00

r456	178	443	4.603000e+00
c457	443	0	4.603e-14
r458	443	444	4.603000e+00
c459	444	0	4.603e-14
r460	444	180	4.603000e+00

r461	178	445	4.605000e+00
c462	445	0	4.605e-14
r463	445	446	4.605000e+00
c464	446	0	4.605e-14
r465	446	181	4.605000e+00

r466	179	447	2.042000e+00
c467	447	0	2.042e-14
r468	447	448	2.042000e+00
c469	448	0	2.042e-14
r470	448	182	2.042000e+00

r471	179	449	2.043000e+00
c472	449	0	2.043e-14
r473	449	450	2.043000e+00
c474	450	0	2.043e-14
r475	450	183	2.043000e+00

r476	180	451	3.408000e+00
c477	451	0	3.408e-14
r478	451	452	3.408000e+00
c479	452	0	3.408e-14
r480	452	75	3.408000e+00

* port 75 - load 3.900000e-02

r481	180	453	3.410000e+00
c482	453	0	3.41e-14
r483	453	454	3.410000e+00
c484	454	0	3.41e-14
r485	454	68	3.410000e+00

* port 68 - load 3.000000e-02

r486	181	455	8.470000e-01
c487	455	0	8.47e-15
r488	455	456	8.470000e-01
c489	456	0	8.47e-15
r490	456	64	8.470000e-01

* port 64 - load 3.000000e-02

r491	181	457	8.480000e-01
c492	457	0	8.48e-15
r493	457	458	8.480000e-01
c494	458	0	8.48e-15
r495	458	62	8.480000e-01

* port 62 - load 5.000000e-02

r496	182	459	1.493000e+00
c497	459	0	1.493e-14
r498	459	460	1.493000e+00
c499	460	0	1.493e-14
r500	460	71	1.493000e+00

* port 71 - load 3.400000e-02

r501	182	461	1.492000e+00
c502	461	0	1.492e-14
r503	461	462	1.492000e+00
c504	462	0	1.492e-14
r505	462	58	1.492000e+00

* port 58 - load 3.200000e-02

r506	183	463	2.032000e+00
c507	463	0	2.032e-14
r508	463	464	2.032000e+00
c509	464	0	2.032e-14
r510	464	60	2.032000e+00

* port 60 - load 6.700000e-02

r511	183	465	2.031000e+00
c512	465	0	2.031e-14
r513	465	466	2.031000e+00
c514	466	0	2.031e-14
r515	466	74	2.031000e+00

* port 74 - load 3.800000e-02

r516	170	467	5.612000e+00
c517	467	0	5.612e-14
r518	467	468	5.612000e+00
c519	468	0	5.612e-14
r520	468	184	5.612000e+00

r521	170	469	5.613000e+00
c522	469	0	5.613e-14
r523	469	470	5.613000e+00
c524	470	0	5.613e-14
r525	470	185	5.613000e+00

r526	184	471	3.829000e+00
c527	471	0	3.829e-14
r528	471	472	3.829000e+00
c529	472	0	3.829e-14
r530	472	186	3.829000e+00

r531	184	473	3.829000e+00
c532	473	0	3.829e-14
r533	473	474	3.829000e+00
c534	474	0	3.829e-14
r535	474	187	3.829000e+00

r536	185	475	5.874000e+00
c537	475	0	5.874e-14
r538	475	476	5.874000e+00
c539	476	0	5.874e-14
r540	476	188	5.874000e+00

r541	185	477	5.874000e+00
c542	477	0	5.874e-14
r543	477	478	5.874000e+00
c544	478	0	5.874e-14
r545	478	189	5.874000e+00

r546	186	479	6.156000e+00
c547	479	0	6.156e-14
r548	479	480	6.156000e+00
c549	480	0	6.156e-14
r550	480	52	6.156000e+00

* port 52 - load 7.400000e-02

r551	186	481	6.157000e+00
c552	481	0	6.157e-14
r553	481	482	6.157000e+00
c554	482	0	6.157e-14
r555	482	66	6.157000e+00

* port 66 - load 5.100000e-02

r556	187	483	3.698000e+00
c557	483	0	3.698e-14
r558	483	484	3.698000e+00
c559	484	0	3.698e-14
r560	484	69	3.698000e+00

* port 69 - load 7.200000e-02

r561	187	485	3.699000e+00
c562	485	0	3.699e-14
r563	485	486	3.699000e+00
c564	486	0	3.699e-14
r565	486	63	3.699000e+00

* port 63 - load 6.900000e-02

r566	188	487	6.282000e+00
c567	487	0	6.282e-14
r568	487	488	6.282000e+00
c569	488	0	6.282e-14
r570	488	2	6.282000e+00

* port 2 - load 3.500000e-02

r571	188	489	6.284000e+00
c572	489	0	6.284e-14
r573	489	490	6.284000e+00
c574	490	0	6.284e-14
r575	490	7	6.284000e+00

* port 7 - load 7.200000e-02

r576	189	491	1.408000e+00
c577	491	0	1.408e-14
r578	491	492	1.408000e+00
c579	492	0	1.408e-14
r580	492	9	1.408000e+00

* port 9 - load 4.500000e-02

r581	189	493	1.409000e+00
c582	493	0	1.409e-14
r583	493	494	1.409000e+00
c584	494	0	1.409e-14
r585	494	3	1.409000e+00

* port 3 - load 5.300000e-02

r586	171	495	4.702000e+00
c587	495	0	4.702e-14
r588	495	496	4.702000e+00
c589	496	0	4.702e-14
r590	496	190	4.702000e+00

r591	171	497	4.703000e+00
c592	497	0	4.703e-14
r593	497	498	4.703000e+00
c594	498	0	4.703e-14
r595	498	191	4.703000e+00

r596	190	499	3.461000e+00
c597	499	0	3.461e-14
r598	499	500	3.461000e+00
c599	500	0	3.461e-14
r600	500	192	3.461000e+00

r601	190	501	3.461000e+00
c602	501	0	3.461e-14
r603	501	502	3.461000e+00
c604	502	0	3.461e-14
r605	502	193	3.461000e+00

r606	191	503	4.176000e+00
c607	503	0	4.176e-14
r608	503	504	4.176000e+00
c609	504	0	4.176e-14
r610	504	194	4.176000e+00

r611	191	505	4.176000e+00
c612	505	0	4.176e-14
r613	505	506	4.176000e+00
c614	506	0	4.176e-14
r615	506	195	4.176000e+00

r616	192	507	2.185000e+00
c617	507	0	2.185e-14
r618	507	508	2.185000e+00
c619	508	0	2.185e-14
r620	508	61	2.185000e+00

* port 61 - load 6.600000e-02

r621	192	509	2.187000e+00
c622	509	0	2.187e-14
r623	509	510	2.187000e+00
c624	510	0	2.187e-14
r625	510	73	2.187000e+00

* port 73 - load 4.600000e-02

r626	193	511	2.125000e+00
c627	511	0	2.125e-14
r628	511	512	2.125000e+00
c629	512	0	2.125e-14
r630	512	59	2.125000e+00

* port 59 - load 7.400000e-02

r631	193	513	2.125000e+00
c632	513	0	2.125e-14
r633	513	514	2.125000e+00
c634	514	0	2.125e-14
r635	514	70	2.125000e+00

* port 70 - load 6.600000e-02

r636	194	515	2.596000e+00
c637	515	0	2.596e-14
r638	515	516	2.596000e+00
c639	516	0	2.596e-14
r640	516	5	2.596000e+00

* port 5 - load 4.500000e-02

r641	194	517	2.596000e+00
c642	517	0	2.596e-14
r643	517	518	2.596000e+00
c644	518	0	2.596e-14
r645	518	4	2.596000e+00

* port 4 - load 3.400000e-02

r646	195	519	2.455000e+00
c647	519	0	2.455e-14
r648	519	520	2.455000e+00
c649	520	0	2.455e-14
r650	520	72	2.455000e+00

* port 72 - load 8.000000e-02

r651	195	521	2.456000e+00
c652	521	0	2.456e-14
r653	521	522	2.456000e+00
c654	522	0	2.456e-14
r655	522	8	2.456000e+00

* port 8 - load 4.300000e-02

r656	134	523	7.103000e+00
c657	523	0	7.103e-14
r658	523	524	7.103000e+00
c659	524	0	7.103e-14
r660	524	196	7.103000e+00

r661	134	525	7.102000e+00
c662	525	0	7.102e-14
r663	525	526	7.102000e+00
c664	526	0	7.102e-14
r665	526	197	7.102000e+00

r666	196	527	6.917000e+00
c667	527	0	6.917e-14
r668	527	528	6.917000e+00
c669	528	0	6.917e-14
r670	528	198	6.917000e+00

r671	196	529	6.915000e+00
c672	529	0	6.915e-14
r673	529	530	6.915000e+00
c674	530	0	6.915e-14
r675	530	199	6.915000e+00

r676	197	531	5.706000e+00
c677	531	0	5.706e-14
r678	531	532	5.706000e+00
c679	532	0	5.706e-14
r680	532	200	5.706000e+00

r681	197	533	5.705000e+00
c682	533	0	5.705e-14
r683	533	534	5.705000e+00
c684	534	0	5.705e-14
r685	534	201	5.705000e+00

r686	198	535	5.489000e+00
c687	535	0	5.489e-14
r688	535	536	5.489000e+00
c689	536	0	5.489e-14
r690	536	202	5.489000e+00

r691	198	537	5.490000e+00
c692	537	0	5.49e-14
r693	537	538	5.490000e+00
c694	538	0	5.49e-14
r695	538	203	5.490000e+00

r696	202	539	5.459000e+00
c697	539	0	5.459e-14
r698	539	540	5.459000e+00
c699	540	0	5.459e-14
r700	540	204	5.459000e+00

r701	202	541	5.458000e+00
c702	541	0	5.458e-14
r703	541	542	5.458000e+00
c704	542	0	5.458e-14
r705	542	205	5.458000e+00

r706	203	543	2.907000e+00
c707	543	0	2.907e-14
r708	543	544	2.907000e+00
c709	544	0	2.907e-14
r710	544	206	2.907000e+00

r711	203	545	2.907000e+00
c712	545	0	2.907e-14
r713	545	546	2.907000e+00
c714	546	0	2.907e-14
r715	546	207	2.907000e+00

r716	204	547	1.660000e+00
c717	547	0	1.66e-14
r718	547	548	1.660000e+00
c719	548	0	1.66e-14
r720	548	121	1.660000e+00

* port 121 - load 7.400000e-02

r721	204	549	1.661000e+00
c722	549	0	1.661e-14
r723	549	550	1.661000e+00
c724	550	0	1.661e-14
r725	550	128	1.661000e+00

* port 128 - load 3.200000e-02

r726	205	551	2.484000e+00
c727	551	0	2.484e-14
r728	551	552	2.484000e+00
c729	552	0	2.484e-14
r730	552	127	2.484000e+00

* port 127 - load 6.700000e-02

r731	205	553	2.484000e+00
c732	553	0	2.484e-14
r733	553	554	2.484000e+00
c734	554	0	2.484e-14
r735	554	122	2.484000e+00

* port 122 - load 3.200000e-02

r736	206	555	2.927000e+00
c737	555	0	2.927e-14
r738	555	556	2.927000e+00
c739	556	0	2.927e-14
r740	556	120	2.927000e+00

* port 120 - load 6.400000e-02

r741	206	557	2.928000e+00
c742	557	0	2.928e-14
r743	557	558	2.928000e+00
c744	558	0	2.928e-14
r745	558	124	2.928000e+00

* port 124 - load 3.300000e-02

r746	207	559	9.940000e-01
c747	559	0	9.94e-15
r748	559	560	9.940000e-01
c749	560	0	9.94e-15
r750	560	106	9.940000e-01

* port 106 - load 3.400000e-02

r751	207	561	9.930000e-01
c752	561	0	9.93e-15
r753	561	562	9.930000e-01
c754	562	0	9.93e-15
r755	562	93	9.930000e-01

* port 93 - load 7.800000e-02

r756	199	563	5.441000e+00
c757	563	0	5.441e-14
r758	563	564	5.441000e+00
c759	564	0	5.441e-14
r760	564	208	5.441000e+00

r761	199	565	5.441000e+00
c762	565	0	5.441e-14
r763	565	566	5.441000e+00
c764	566	0	5.441e-14
r765	566	209	5.441000e+00

r766	208	567	1.174000e+00
c767	567	0	1.174e-14
r768	567	568	1.174000e+00
c769	568	0	1.174e-14
r770	568	210	1.174000e+00

r771	208	569	1.173000e+00
c772	569	0	1.173e-14
r773	569	570	1.173000e+00
c774	570	0	1.173e-14
r775	570	211	1.173000e+00

r776	209	571	3.888000e+00
c777	571	0	3.888e-14
r778	571	572	3.888000e+00
c779	572	0	3.888e-14
r780	572	212	3.888000e+00

r781	209	573	3.890000e+00
c782	573	0	3.89e-14
r783	573	574	3.890000e+00
c784	574	0	3.89e-14
r785	574	213	3.890000e+00

r786	210	575	2.552000e+00
c787	575	0	2.552e-14
r788	575	576	2.552000e+00
c789	576	0	2.552e-14
r790	576	25	2.552000e+00

* port 25 - load 3.700000e-02

r791	210	577	2.552000e+00
c792	577	0	2.552e-14
r793	577	578	2.552000e+00
c794	578	0	2.552e-14
r795	578	105	2.552000e+00

* port 105 - load 5.000000e-02

r796	211	579	3.088000e+00
c797	579	0	3.088e-14
r798	579	580	3.088000e+00
c799	580	0	3.088e-14
r800	580	90	3.088000e+00

* port 90 - load 6.000000e-02

r801	211	581	3.088000e+00
c802	581	0	3.088e-14
r803	581	582	3.088000e+00
c804	582	0	3.088e-14
r805	582	30	3.088000e+00

* port 30 - load 3.200000e-02

r806	212	583	5.050000e+00
c807	583	0	5.05e-14
r808	583	584	5.050000e+00
c809	584	0	5.05e-14
r810	584	92	5.050000e+00

* port 92 - load 4.100000e-02

r811	212	585	5.050000e+00
c812	585	0	5.05e-14
r813	585	586	5.050000e+00
c814	586	0	5.05e-14
r815	586	104	5.050000e+00

* port 104 - load 6.600000e-02

r816	213	587	4.330000e+00
c817	587	0	4.33e-14
r818	587	588	4.330000e+00
c819	588	0	4.33e-14
r820	588	31	4.330000e+00

* port 31 - load 6.000000e-02

r821	213	589	4.330000e+00
c822	589	0	4.33e-14
r823	589	590	4.330000e+00
c824	590	0	4.33e-14
r825	590	125	4.330000e+00

* port 125 - load 6.400000e-02

r826	200	591	5.099000e+00
c827	591	0	5.099e-14
r828	591	592	5.099000e+00
c829	592	0	5.099e-14
r830	592	214	5.099000e+00

r831	200	593	5.099000e+00
c832	593	0	5.099e-14
r833	593	594	5.099000e+00
c834	594	0	5.099e-14
r835	594	215	5.099000e+00

r836	214	595	4.677000e+00
c837	595	0	4.677e-14
r838	595	596	4.677000e+00
c839	596	0	4.677e-14
r840	596	216	4.677000e+00

r841	214	597	4.679000e+00
c842	597	0	4.679e-14
r843	597	598	4.679000e+00
c844	598	0	4.679e-14
r845	598	217	4.679000e+00

r846	215	599	3.842000e+00
c847	599	0	3.842e-14
r848	599	600	3.842000e+00
c849	600	0	3.842e-14
r850	600	218	3.842000e+00

r851	215	601	3.844000e+00
c852	601	0	3.844e-14
r853	601	602	3.844000e+00
c854	602	0	3.844e-14
r855	602	219	3.844000e+00

r856	216	603	3.154000e+00
c857	603	0	3.154e-14
r858	603	604	3.154000e+00
c859	604	0	3.154e-14
r860	604	119	3.154000e+00

* port 119 - load 5.800000e-02

r861	216	605	3.155000e+00
c862	605	0	3.155e-14
r863	605	606	3.155000e+00
c864	606	0	3.155e-14
r865	606	123	3.155000e+00

* port 123 - load 5.400000e-02

r866	217	607	2.183000e+00
c867	607	0	2.183e-14
r868	607	608	2.183000e+00
c869	608	0	2.183e-14
r870	608	118	2.183000e+00

* port 118 - load 7.600000e-02

r871	217	609	2.183000e+00
c872	609	0	2.183e-14
r873	609	610	2.183000e+00
c874	610	0	2.183e-14
r875	610	115	2.183000e+00

* port 115 - load 3.600000e-02

r876	218	611	2.651000e+00
c877	611	0	2.651e-14
r878	611	612	2.651000e+00
c879	612	0	2.651e-14
r880	612	112	2.651000e+00

* port 112 - load 3.300000e-02

r881	218	613	2.652000e+00
c882	613	0	2.652e-14
r883	613	614	2.652000e+00
c884	614	0	2.652e-14
r885	614	113	2.652000e+00

* port 113 - load 4.400000e-02

r886	219	615	3.126000e+00
c887	615	0	3.126e-14
r888	615	616	3.126000e+00
c889	616	0	3.126e-14
r890	616	114	3.126000e+00

* port 114 - load 5.000000e-02

r891	219	617	3.127000e+00
c892	617	0	3.127e-14
r893	617	618	3.127000e+00
c894	618	0	3.127e-14
r895	618	111	3.127000e+00

* port 111 - load 6.600000e-02

r896	201	619	2.686000e+00
c897	619	0	2.686e-14
r898	619	620	2.686000e+00
c899	620	0	2.686e-14
r900	620	220	2.686000e+00

r901	201	621	2.686000e+00
c902	621	0	2.686e-14
r903	621	622	2.686000e+00
c904	622	0	2.686e-14
r905	622	221	2.686000e+00

r906	220	623	4.025000e+00
c907	623	0	4.025e-14
r908	623	624	4.025000e+00
c909	624	0	4.025e-14
r910	624	222	4.025000e+00

r911	220	625	4.025000e+00
c912	625	0	4.025e-14
r913	625	626	4.025000e+00
c914	626	0	4.025e-14
r915	626	223	4.025000e+00

r916	221	627	3.096000e+00
c917	627	0	3.096e-14
r918	627	628	3.096000e+00
c919	628	0	3.096e-14
r920	628	224	3.096000e+00

r921	221	629	3.098000e+00
c922	629	0	3.098e-14
r923	629	630	3.098000e+00
c924	630	0	3.098e-14
r925	630	225	3.098000e+00

r926	222	631	3.131000e+00
c927	631	0	3.131e-14
r928	631	632	3.131000e+00
c929	632	0	3.131e-14
r930	632	126	3.131000e+00

* port 126 - load 4.000000e-02

r931	222	633	3.132000e+00
c932	633	0	3.132e-14
r933	633	634	3.132000e+00
c934	634	0	3.132e-14
r935	634	116	3.132000e+00

* port 116 - load 4.800000e-02

r936	223	635	1.279000e+00
c937	635	0	1.279e-14
r938	635	636	1.279000e+00
c939	636	0	1.279e-14
r940	636	103	1.279000e+00

* port 103 - load 7.000000e-02

r941	223	637	1.279000e+00
c942	637	0	1.279e-14
r943	637	638	1.279000e+00
c944	638	0	1.279e-14
r945	638	94	1.279000e+00

* port 94 - load 7.200000e-02

r946	224	639	3.697000e+00
c947	639	0	3.697e-14
r948	639	640	3.697000e+00
c949	640	0	3.697e-14
r950	640	110	3.697000e+00

* port 110 - load 7.300000e-02

r951	224	641	3.696000e+00
c952	641	0	3.696e-14
r953	641	642	3.696000e+00
c954	642	0	3.696e-14
r955	642	117	3.696000e+00

* port 117 - load 4.000000e-02

r956	225	643	3.328000e+00
c957	643	0	3.328e-14
r958	643	644	3.328000e+00
c959	644	0	3.328e-14
r960	644	107	3.328000e+00

* port 107 - load 5.100000e-02

r961	225	645	3.329000e+00
c962	645	0	3.329e-14
r963	645	646	3.329000e+00
c964	646	0	3.329e-14
r965	646	100	3.329000e+00

* port 100 - load 6.500000e-02

r966	135	647	1.138200e+01
c967	647	0	1.1382e-13
r968	647	648	1.138200e+01
c969	648	0	1.1382e-13
r970	648	226	1.138200e+01

r971	135	649	1.138100e+01
c972	649	0	1.1381e-13
r973	649	650	1.138100e+01
c974	650	0	1.1381e-13
r975	650	227	1.138100e+01

r976	226	651	1.297900e+01
c977	651	0	1.2979e-13
r978	651	652	1.297900e+01
c979	652	0	1.2979e-13
r980	652	228	1.297900e+01

r981	226	653	1.298000e+01
c982	653	0	1.298e-13
r983	653	654	1.298000e+01
c984	654	0	1.298e-13
r985	654	229	1.298000e+01

r986	227	655	8.838000e+00
c987	655	0	8.838e-14
r988	655	656	8.838000e+00
c989	656	0	8.838e-14
r990	656	230	8.838000e+00

r991	227	657	8.838000e+00
c992	657	0	8.838e-14
r993	657	658	8.838000e+00
c994	658	0	8.838e-14
r995	658	231	8.838000e+00

r996	228	659	3.403000e+00
c997	659	0	3.403e-14
r998	659	660	3.403000e+00
c999	660	0	3.403e-14
r1000	660	232	3.403000e+00

r1001	228	661	3.403000e+00
c1002	661	0	3.403e-14
r1003	661	662	3.403000e+00
c1004	662	0	3.403e-14
r1005	662	233	3.403000e+00

r1006	232	663	4.676000e+00
c1007	663	0	4.676e-14
r1008	663	664	4.676000e+00
c1009	664	0	4.676e-14
r1010	664	234	4.676000e+00

r1011	232	665	4.677000e+00
c1012	665	0	4.677e-14
r1013	665	666	4.677000e+00
c1014	666	0	4.677e-14
r1015	666	235	4.677000e+00

r1016	233	667	1.672000e+00
c1017	667	0	1.672e-14
r1018	667	668	1.672000e+00
c1019	668	0	1.672e-14
r1020	668	236	1.672000e+00

r1021	233	669	1.672000e+00
c1022	669	0	1.672e-14
r1023	669	670	1.672000e+00
c1024	670	0	1.672e-14
r1025	670	237	1.672000e+00

r1026	234	671	1.088000e+00
c1027	671	0	1.088e-14
r1028	671	672	1.088000e+00
c1029	672	0	1.088e-14
r1030	672	91	1.088000e+00

* port 91 - load 7.600000e-02

r1031	234	673	1.089000e+00
c1032	673	0	1.089e-14
r1033	673	674	1.089000e+00
c1034	674	0	1.089e-14
r1035	674	29	1.089000e+00

* port 29 - load 6.500000e-02

r1036	235	675	8.710000e-01
c1037	675	0	8.71e-15
r1038	675	676	8.710000e-01
c1039	676	0	8.71e-15
r1040	676	35	8.710000e-01

* port 35 - load 7.300000e-02

r1041	235	677	8.700000e-01
c1042	677	0	8.7e-15
r1043	677	678	8.700000e-01
c1044	678	0	8.7e-15
r1045	678	28	8.700000e-01

* port 28 - load 4.600000e-02

r1046	236	679	2.186000e+00
c1047	679	0	2.186e-14
r1048	679	680	2.186000e+00
c1049	680	0	2.186e-14
r1050	680	34	2.186000e+00

* port 34 - load 7.100000e-02

r1051	236	681	2.186000e+00
c1052	681	0	2.186e-14
r1053	681	682	2.186000e+00
c1054	682	0	2.186e-14
r1055	682	33	2.186000e+00

* port 33 - load 4.000000e-02

r1056	237	683	2.530000e+00
c1057	683	0	2.53e-14
r1058	683	684	2.530000e+00
c1059	684	0	2.53e-14
r1060	684	24	2.530000e+00

* port 24 - load 6.800000e-02

r1061	237	685	2.530000e+00
c1062	685	0	2.53e-14
r1063	685	686	2.530000e+00
c1064	686	0	2.53e-14
r1065	686	23	2.530000e+00

* port 23 - load 6.500000e-02

r1066	229	687	1.468300e+01
c1067	687	0	1.4683e-13
r1068	687	688	1.468300e+01
c1069	688	0	1.4683e-13
r1070	688	238	1.468300e+01

r1071	229	689	1.468300e+01
c1072	689	0	1.4683e-13
r1073	689	690	1.468300e+01
c1074	690	0	1.4683e-13
r1075	690	239	1.468300e+01

r1076	238	691	3.556000e+00
c1077	691	0	3.556e-14
r1078	691	692	3.556000e+00
c1079	692	0	3.556e-14
r1080	692	240	3.556000e+00

r1081	238	693	3.556000e+00
c1082	693	0	3.556e-14
r1083	693	694	3.556000e+00
c1084	694	0	3.556e-14
r1085	694	241	3.556000e+00

r1086	239	695	6.675000e+00
c1087	695	0	6.675e-14
r1088	695	696	6.675000e+00
c1089	696	0	6.675e-14
r1090	696	242	6.675000e+00

r1091	239	697	6.675000e+00
c1092	697	0	6.675e-14
r1093	697	698	6.675000e+00
c1094	698	0	6.675e-14
r1095	698	243	6.675000e+00

r1096	240	699	3.164000e+00
c1097	699	0	3.164e-14
r1098	699	700	3.164000e+00
c1099	700	0	3.164e-14
r1100	700	11	3.164000e+00

* port 11 - load 3.300000e-02

r1101	240	701	3.165000e+00
c1102	701	0	3.165e-14
r1103	701	702	3.165000e+00
c1104	702	0	3.165e-14
r1105	702	12	3.165000e+00

* port 12 - load 3.200000e-02

r1106	241	703	4.208000e+00
c1107	703	0	4.208e-14
r1108	703	704	4.208000e+00
c1109	704	0	4.208e-14
r1110	704	6	4.208000e+00

* port 6 - load 7.000000e-02

r1111	241	705	4.209000e+00
c1112	705	0	4.209e-14
r1113	705	706	4.209000e+00
c1114	706	0	4.209e-14
r1115	706	10	4.209000e+00

* port 10 - load 4.300000e-02

r1116	242	707	6.984000e+00
c1117	707	0	6.984e-14
r1118	707	708	6.984000e+00
c1119	708	0	6.984e-14
r1120	708	32	6.984000e+00

* port 32 - load 7.800000e-02

r1121	242	709	6.985000e+00
c1122	709	0	6.985e-14
r1123	709	710	6.985000e+00
c1124	710	0	6.985e-14
r1125	710	18	6.985000e+00

* port 18 - load 3.700000e-02

r1126	243	711	1.732000e+00
c1127	711	0	1.732e-14
r1128	711	712	1.732000e+00
c1129	712	0	1.732e-14
r1130	712	15	1.732000e+00

* port 15 - load 4.300000e-02

r1131	243	713	1.733000e+00
c1132	713	0	1.733e-14
r1133	713	714	1.733000e+00
c1134	714	0	1.733e-14
r1135	714	14	1.733000e+00

* port 14 - load 6.700000e-02

r1136	230	715	4.261000e+00
c1137	715	0	4.261e-14
r1138	715	716	4.261000e+00
c1139	716	0	4.261e-14
r1140	716	244	4.261000e+00

r1141	230	717	4.261000e+00
c1142	717	0	4.261e-14
r1143	717	718	4.261000e+00
c1144	718	0	4.261e-14
r1145	718	245	4.261000e+00

r1146	244	719	4.373000e+00
c1147	719	0	4.373e-14
r1148	719	720	4.373000e+00
c1149	720	0	4.373e-14
r1150	720	246	4.373000e+00

r1151	244	721	4.373000e+00
c1152	721	0	4.373e-14
r1153	721	722	4.373000e+00
c1154	722	0	4.373e-14
r1155	722	247	4.373000e+00

r1156	245	723	1.966000e+00
c1157	723	0	1.966e-14
r1158	723	724	1.966000e+00
c1159	724	0	1.966e-14
r1160	724	248	1.966000e+00

r1161	245	725	1.967000e+00
c1162	725	0	1.967e-14
r1163	725	726	1.967000e+00
c1164	726	0	1.967e-14
r1165	726	249	1.967000e+00

r1166	246	727	7.760000e-01
c1167	727	0	7.76e-15
r1168	727	728	7.760000e-01
c1169	728	0	7.76e-15
r1170	728	95	7.760000e-01

* port 95 - load 7.500000e-02

r1171	246	729	7.780000e-01
c1172	729	0	7.78e-15
r1173	729	730	7.780000e-01
c1174	730	0	7.78e-15
r1175	730	97	7.780000e-01

* port 97 - load 7.000000e-02

r1176	247	731	4.364000e+00
c1177	731	0	4.364e-14
r1178	731	732	4.364000e+00
c1179	732	0	4.364e-14
r1180	732	101	4.364000e+00

* port 101 - load 5.200000e-02

r1181	247	733	4.365000e+00
c1182	733	0	4.365e-14
r1183	733	734	4.365000e+00
c1184	734	0	4.365e-14
r1185	734	96	4.365000e+00

* port 96 - load 3.300000e-02

r1186	248	735	3.087000e+00
c1187	735	0	3.087e-14
r1188	735	736	3.087000e+00
c1189	736	0	3.087e-14
r1190	736	108	3.087000e+00

* port 108 - load 4.800000e-02

r1191	248	737	3.087000e+00
c1192	737	0	3.087e-14
r1193	737	738	3.087000e+00
c1194	738	0	3.087e-14
r1195	738	109	3.087000e+00

* port 109 - load 6.900000e-02

r1196	249	739	4.194000e+00
c1197	739	0	4.194e-14
r1198	739	740	4.194000e+00
c1199	740	0	4.194e-14
r1200	740	102	4.194000e+00

* port 102 - load 5.400000e-02

r1201	249	741	4.196000e+00
c1202	741	0	4.196e-14
r1203	741	742	4.196000e+00
c1204	742	0	4.196e-14
r1205	742	99	4.196000e+00

* port 99 - load 3.800000e-02

r1206	231	743	6.918000e+00
c1207	743	0	6.918e-14
r1208	743	744	6.918000e+00
c1209	744	0	6.918e-14
r1210	744	250	6.918000e+00

r1211	231	745	6.917000e+00
c1212	745	0	6.917e-14
r1213	745	746	6.917000e+00
c1214	746	0	6.917e-14
r1215	746	251	6.917000e+00

r1216	250	747	7.988000e+00
c1217	747	0	7.988e-14
r1218	747	748	7.988000e+00
c1219	748	0	7.988e-14
r1220	748	252	7.988000e+00

r1221	250	749	7.987000e+00
c1222	749	0	7.987e-14
r1223	749	750	7.987000e+00
c1224	750	0	7.987e-14
r1225	750	253	7.987000e+00

r1226	251	751	6.202000e+00
c1227	751	0	6.202e-14
r1228	751	752	6.202000e+00
c1229	752	0	6.202e-14
r1230	752	254	6.202000e+00

r1231	251	753	6.201000e+00
c1232	753	0	6.201e-14
r1233	753	754	6.201000e+00
c1234	754	0	6.201e-14
r1235	754	255	6.201000e+00

r1236	252	755	1.323000e+00
c1237	755	0	1.323e-14
r1238	755	756	1.323000e+00
c1239	756	0	1.323e-14
r1240	756	22	1.323000e+00

* port 22 - load 4.000000e-02

r1241	252	757	1.323000e+00
c1242	757	0	1.323e-14
r1243	757	758	1.323000e+00
c1244	758	0	1.323e-14
r1245	758	17	1.323000e+00

* port 17 - load 4.000000e-02

r1246	253	759	1.089200e+01
c1247	759	0	1.0892e-13
r1248	759	760	1.089200e+01
c1249	760	0	1.0892e-13
r1250	760	13	1.089200e+01

* port 13 - load 3.100000e-02

r1251	253	761	1.089100e+01
c1252	761	0	1.0891e-13
r1253	761	762	1.089100e+01
c1254	762	0	1.0891e-13
r1255	762	16	1.089100e+01

* port 16 - load 3.500000e-02

r1256	254	763	1.971000e+00
c1257	763	0	1.971e-14
r1258	763	764	1.971000e+00
c1259	764	0	1.971e-14
r1260	764	20	1.971000e+00

* port 20 - load 5.300000e-02

r1261	254	765	1.970000e+00
c1262	765	0	1.97e-14
r1263	765	766	1.970000e+00
c1264	766	0	1.97e-14
r1265	766	98	1.970000e+00

* port 98 - load 3.700000e-02

r1266	255	767	2.388000e+00
c1267	767	0	2.388e-14
r1268	767	768	2.388000e+00
c1269	768	0	2.388e-14
r1270	768	19	2.388000e+00

* port 19 - load 5.500000e-02

r1271	255	769	2.387000e+00
c1272	769	0	2.387e-14
r1273	769	770	2.387000e+00
c1274	770	0	2.387e-14
r1275	770	21	2.387000e+00

* port 21 - load 6.300000e-02

*AC analysis
*.AC 100 1e7 1e9 
.RD PRIMA
*report results
*.PLOTNV 769
*.PLOTNV 41
