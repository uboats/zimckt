* circuit described in the handout
*Vin 101 0 PWL 0 0 5.0e-10 3.0
*Rin 101 102 10
*L1  102 103 1e-7
*R1 103 104 10
*C1 104 0 0.1e-12

R1 101 0 10
R2 101 102 10
*I1 0 102 PWL 0 0 5.0e-10 0.2 1e-9 0.2 1.5e-9 0.1
I1 0 102 SIN 0 0.1 10000 0

*.DC
.TRAN TR 1e-5 1.0e-3
*.TRAN TR 1e-12 2.0e-9
.PLOTNV 101
.PLOTNV 102


*.TRAN TR 1e-12 2.0e-9
*.PLOTNV 104
*.PLOTNV 101
*.PLOTNV 102
*.PLOTNV 103
