* ckt file for parser

* interpret this as a voltage step

Idriver1 1 0 1
r6 4 0 10

* port 256 - load 2.000000e+00

r1	1	2	1
c2  2	0	1e-6
r3	2	3	1
c4	3	0	1e-6
r5	3	4	1
c4	4	0	1e-6

.RD PRIMA
