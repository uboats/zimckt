* circuit described in the handout
*Vin 101 0 PWL 0 0 5.0e-10 3.0
Vin 101 0 SIN 0 0.1 10000 0
*Vin 101 0 PULSE 0.1 2 5e-5 10e-5 5e-5 10e-5 3e-4
VDD 103 0 DC 10

C1 101 102 10e-6
Rg1 102 0 2000
R1 103 102 8000
R3 103 104 150000
Rl 105 0 10000
Cl 104 105 10e-6


M1 104 102 0 n 10e-6 0.35e-6 2
.MODEL 2 VT 0.83 MU 1.5e-1 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14

.TRAN TR 1e-5 1.0e-3

.PLOTNV 101
.PLOTNV 105
*.PLOTNV 103
*.PLOTNV 104
