* ac test

vin 101 0 AC 2
R1 101 102 2
L1 102 0 2.5e-5
L2 102 103 2.5e-6
Rl 103 0 100

*.AC LIN  500 10 1000
.AC DEC 20 10 5000000000
*.PLOTNV 102
.PLOTNV 103